module fifo_3();
endmodule
