module mul_2x2();

endmodule
