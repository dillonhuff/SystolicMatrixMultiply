module inner_product_3();
endmodule
